library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use std.textio.all;

entity sync_ram is
  port (
    clock   : in  std_logic;
    w_en      : in  std_logic;
    address : in  std_logic_vector(31 downto 0);
    datain  : in  std_logic_vector(31 downto 0);
    dataout : out std_logic_vector(31 downto 0)
  );
end entity sync_ram;

architecture RTL of sync_ram is

   type ram_type is array (0 to (2**32)-1) of std_logic_vector(31 downto 0);
   signal ram : ram_type;
   signal read_address : std_logic_vector(31 downto 0);
	signal lida : std_logic := '0';
begin

  
  impure function ReadMemFile(FileName : STRING) return ram_type is
  file FileHandle       : TEXT open READ_MODE is FileName;
  variable CurrentLine  : LINE;
  variable TempWord     : bit_vector(31 downto 0);
  variable Result       : ram_type    := (others => (others => '0'));

  RamProc: process(clock) is

  begin
	if lida = '0' then
		for i in 0 to 4095 loop
			 exit when endfile(FileHandle);
			 readline(FileHandle, CurrentLine);
			 read(CurrentLine, TempWord);
			 Result(i) := to_stdlogicvector(TempWord);
		 end loop;
		 lida = '1';
	end if 
  
    if rising_edge(clock) then
      if w_en = '1' then
        ram(to_integer(unsigned(address))) <= datain;
      end if;
      read_address <= address;
    end if;
  end process RamProc;

  dataout <= ram(to_integer(unsigned(read_address)));

end architecture RTL;


