library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alu is 
    port (
        in_1, in_2: std_logic_vector(31 downto 0);
        alu_control_funct: in std_logic_vector(3 downto 0);
        zero: out std_logic;
        alu_result: out std_logic_vector(31 downto 0)
    );
end alu;

architecture beh of alu is
begin
    process(alu_control_funct, in_1, in_2)
    begin
        case alu_control_funct is
            when "0010" => -- add
                alu_result <= in_1 + in_2;
            when "0110" => -- subtract
                alu_result <=  in_1 - in_2;
            when "0011" => -- subtract not equal
                alu_result <=  in_1 - in_2;
            when "0000" => -- and
                alu_result <= in_1 and in_2;
            when "0001" => -- or
                alu_result <= in_1 or in_2;
            when "0111" => -- set on less than
                if in_1 < in_2 then
                    alu_result <= "00000000000000000000000000000001";
                else
                    alu_result <= "00000000000000000000000000000000";
                end if;
            when others =>
                alu_result <= (others => 'X');
        end case;

        if alu_control_funct = "0011" then -- subtract not equal
            if in_1 = in_2 then
                zero <= '0';
            else
                zero <= '1';
            end if;
        else
            if in_1 = in_2 then
                zero <= '1';
            else
                zero <= '0';
            end if;
        end if;
    end process;
end beh;
