library IEEE;
use IEEE.std_logic_1164.all;

entity extensor_8to32 is
    port (
        data_in: in std_logic_vector(7 downto 0);
        data_out: out std_logic_vector(31 downto 0)
    );
end extensor_8to32;

architecture beh of extensor_8to32 is
begin
    process(data_in)
    begin
        data_out <= (others => '0');
        data_out(7 downto 0) <= data_in;
    end process;
end beh;
